q1.1
v 1 0 dc pulse(0 1 0 0 0 100u)
r 2 0 1k
c 1 2 10n
.tran 0.1us 100us
.control
run
plot v(2)/1000
hardcopy q1_1 v(2)/1000
.endc
.end
