*Ids-Vds and Ids-Vgs of a n-MOSFET
.include tsmc.txt
M1 2 1 0 0 CMOSN W=10u
VDD 2 0 DC 5v
VGG 1 0 DC 3.85V

*defining the run-time control functions
.dc VGG 0 5 0.05 
*VDD 0 5 5
*.dc VDD 0 10 0.05
.control

run
*plotting input and output voltages
plot -I(vdd)
*plot deriv(-I(vdd))
*plot I(vgg) vs v(1)
hardcopy q1 -I(vdd)
.endc
.end
