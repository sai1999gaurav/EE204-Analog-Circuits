*Ids-Vds and Ids-Vgs of a n-MOSFET
.include tsmc.txt
M1 2 1 0 0 CMOSN W=10u
VDD 3 0 dc 15v
Vgg 4 0 dc 2.1v
Rd 2 3 19k
Vin 1 4 ac sin(0 100m 1k 0 0)
.tran 0.02m 10m
.control
run
plot (v(1)-v(4)),  v(2)-4
hardcopy q1 (v(1)-v(4)),  v(2)-4
.endc
.end 
