q1.1
v1 1 0 ac 1
r1 1 2 1k
c1 2 0 10n
v2 3 0 ac 1
r2 3 4 1k
c2 4 5 10n
l2 5 0 1m
v3 6 0 ac 1
r3 6 7 1k
l3 7 0 1m
.ac lin 1000 0 5000k
.control
run
plot cph(v(1)/i(v1)), cph(v(3)/i(v2)), cph(v(6)/i(v3))
hardcopy q3_1 cph(v(1)/i(v1)), cph(v(3)/i(v2)), cph(v(6)/i(v3))
.endc
.end
