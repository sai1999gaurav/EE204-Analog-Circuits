*wein
.include ua741.txt
X1 2 1 3 4 15 ua741
Vdd 3 0 dc 5v
vss 4 0 dc -5v
vin 7 0 sin(0 1n 100k 0 1u)
r1 1 7 1k
r2 1 15 2k
r3 15 6 10k
c3 6 2 16n
r4 2 0 10k
c4 2 0 16n

.tran 0.01ms 5ms
.control
run
plot V(15)
.endc
.end
