q1.1
v 1 0 sin(0 1 100k -2.5u 1e-10)
r 2 0 1k
c 1 2 10n
.tran 0.001us 100us
.control
run
plot v(1)
plot v(2)/1000
hardcopy q2_1 v(2)/1000
.endc
.end

